//  Class: alu_vseqr
//
class alu_vseqr extends uvm_component;
  `uvm_component_utils(alu_vseqr)


  //  Group: Components


  //  Group: Variables


  //  Group: Functions

  //  Constructor: new
  function new(string name = "alu_vseqr", uvm_component parent);
    super.new(name, parent);
  endfunction : new


endclass : alu_vseqr
