//==============================================================================
// Project: AXI-Stream VIP
//==============================================================================
// Filename: spi_txn.sv
// Description: This file comprises the packet item for AXIS VIP.
//    - This time holds all the data to be transferred in an packet transaction.
//    - It also has a protected transfer queue, which holds the items for
//      independent transfers. These are received by the main driver for the 
//      transfer.
//==============================================================================

//  Class: axis_packet
//
class axis_packet extends uvm_sequence_item;
    // `uvm_object_utils(axis_packet)

  //  Group: Variables

  /* p_data:
      - packet data. should be sent in transfers by transmitter driver.
      - keep and strb are generated as well to allow full randomization,
        when necessary.
  */
  rand bit [TDATA_WIDTH-1:0] p_data[$];
  rand bit [(TDATA_WIDTH/8)-1:0] p_keep[$];
  rand bit [(TDATA_WIDTH/8)-1:0] p_strb[$];


  /* size:
      - number of transfers in this packet.
  */
  rand int size;

  /* delay:
      - Holds a delay to be applied prior to sending this item.
      - This delay is an integer and represents a number of clock cycles.
      NOTE: perhaps delay should be associated with the trasfer and not with
            the packet. If that's the case, it should likely be a queue of delays
            not a single value.
  */
  rand int unsigned delay;

  /* timestamp:
      - Holds the time in which the item was received.
  */
  time timestamps[$];


  /* transfers:
      - holds all transfers collected by the monitor, or generated by the
      transfer2packet converter.
  */
  protected axis_transfer transfers[];


  //  Group: Constraints
  constraint size_c {
    solve size before p_data;

    soft size inside {[1 : 100]};
    p_data.size() == size;
  }

  constraint delay_c {soft delay inside {[0 : 1000]};}

  // Group: Functions
  /* Function: packet2transfer
      Description:
      - Converts the current packet into transfer and builds
      the transfer dynamic array.
  */
  virtual function void packet2transfer();
    string report_id = $sformatf("%s.packet2trasnfer", this.report_id);

    if (this.p_data.size() == 0)
      `uvm_fatal(report_id, $sformatf(
                 {
                   "The item '%s', type of '%s', currently ",
                   "has no data to be converted into trasnfers. Only call this method ",
                   "if the '%s' is ready to be converted into transfers."
                 },
                 this.get_name(),
                 this.get_type(),
                 this.get_type()
                 ))

    if ((this.timestamps.size() != this.p_data.size()) && (this.timestamps.size() > 0))
      `uvm_fatal(report_id, $sformatf(
                 {
                   "The 'timestamps' queue isn't empty, but ",
                   "its size doesn't match the data queue's. ",
                   "Data size: %0d, Timestamps size: %0d"
                 },
                 this.p_data.size(),
                 this.timestamps.size()
                 ))

    transfers = new[this.p_data.size()];

    foreach (this.p_data[i]) begin
      string transfer_name = $sformatf("transfer_%0d", i);

      transfers[i] = axis_transfer::type_id::create(transfer_name);
      transfers[i].tdata = this.p_data[i];
      transfers[i].tkeep = this.p_keep[i];
      transfers[i].tstrb = this.p_strb[i];

      if (this.timestamps.size() > 0) begin
        transfers[i].timestamp = this.timestamps[i];
        transfers[i].delay = i == 0 ? delay : 0;
        transfers[i].tlast = i == p_data.size() - 1;
      end
    end
  endfunction : packet2transfer


  virtual function get_size;
    get_size = this.beats.size();
  endfunction : get_size

  virtual function axis_transfer get_transfer(int i);
    if (i >= this.beats.size())
      `uvm_fatal(this.report_id, "Transfer cannot be retrieved. Array too small for index")
    get_transfer = this.beats[i];
  endfunction : get_transfer


  //  Constructor: new
  function new(string name = "axis_packet");
    super.new(name);
  endfunction : new

  //  Function: do_copy
  // extern function void do_copy(uvm_object rhs);
  //  Function: do_compare
  // extern function bit do_compare(uvm_object rhs, uvm_comparer comparer);
  //  Function: convert2string
  // extern function string convert2string();
  //  Function: do_print
  // extern function void do_print(uvm_printer printer);
  //  Function: do_record
  // extern function void do_record(uvm_recorder recorder);
  //  Function: do_pack
  // extern function void do_pack();
  //  Function: do_unpack
  // extern function void do_unpack();

endclass : axis_packet


/*----------------------------------------------------------------------------*/
/*  Constraints                                                               */
/*----------------------------------------------------------------------------*/




/*----------------------------------------------------------------------------*/
/*  Functions                                                                 */
/*----------------------------------------------------------------------------*/

