
//  Class: axis_packet
//
class axis_packet extends uvm_sequence_item;
  `uvm_object_utils(axis_packet)

  //  Group: Variables

  /* p_data:
      - packet data. should be sent in transfers by transmitter driver.
  */
  rand byte p_data[$];


  /* size:
      - number of transfers in this packet.
  */
  rand int size;

  /* delay:
      - Holds a delay to be applied prior to sending this item.
      - This delay is an integer and represents a number of clock cycles.
  */
  rand int unsigned delay;

  /* timestamp:
      - Holds the time in which the item was received.
  */
  time timestamps[$];


  /* transfers:
      - holds all transfers collected by the monitor, or generated by the
      transfer2packet converter.
  */
  protected axis_transfer transfers[];


  //  Group: Constraints


  //  Group: Functions
  /* Function: packet2transfer

      Description:
      - Converts the current packet into transfer and builds
      the transfer dynamic array.
  */
  virtual function void packet2transfer();
      string report_id = $sformatf("%s.packet2trasnfer", this.report_id);

      if (this.data.size() == 0)
      `uvm_fatal(report_id, $sformatf({"The item '%s', type of '%s', currently ",
                  "has no data to be converted into trasnfers. Only call this method ",
                  "if the '%s' is ready to be converted into transfers."},
                  this.get_name(), this.get_type(), this.get_type()))

      if ((this.timestamps.size() != this.data.size()) &&
          (this.timestamps.size() > 0))
      `uvm_fatal(report_id, $sformatf({"The 'timestamps' queue isn't empty, but ",
                  "its size doesn't match the data queue's. ",
                  "Data size: %0d, Timestamps size: %0d"}, this.data.size(),
                  this.timestamps.size()))

      transfers = new[this.data.size()];

      foreach(this.data[i]) begin
          string transfer_name = $sformatf("transfer_%0d", i);

          transfers[i] = axis_transfer::type_id::create(transfer_name);
          transfers[i].data = this.data[i];

          if (this.timestamps.size() > 0) begin
              transfers[i].timestamp = this.timestamps[i];
              transfers[i].delay = i == 0 ? delay : 0;
              transfers[i].tlast = i == data.size() - 1;
          end

      end
  endfunction : txn2beat_converter



  //  Constructor: new
  function new(string name = "axis_packet");
      super.new(name);
  endfunction: new

  //  Function: do_copy
  // extern function void do_copy(uvm_object rhs);
  //  Function: do_compare
  // extern function bit do_compare(uvm_object rhs, uvm_comparer comparer);
  //  Function: convert2string
  // extern function string convert2string();
  //  Function: do_print
  // extern function void do_print(uvm_printer printer);
  //  Function: do_record
  // extern function void do_record(uvm_recorder recorder);
  //  Function: do_pack
  // extern function void do_pack();
  //  Function: do_unpack
  // extern function void do_unpack();

endclass: axis_packet


/*----------------------------------------------------------------------------*/
/*  Constraints                                                               */
/*----------------------------------------------------------------------------*/




/*----------------------------------------------------------------------------*/
/*  Functions                                                                 */
/*----------------------------------------------------------------------------*/

