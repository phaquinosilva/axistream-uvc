//==============================================================================
// Project: AXI-Stream VIP
//==============================================================================
// Filename: axis_monitor.sv
// Description: This file comprises the monitor of the AXI-Stream VIP.
//==============================================================================
`ifndef axis_monitor__sv
`define axis_monitor__sv 


class axis_monitor extends uvm_monitor;
  `uvm_component_utils(axis_monitor)

  //  Group: Components
  vif_t vif;

  //  Group: Variables
  uvm_analysis_port #(axis_transfer) transfer_ap;
  axis_config m_cfg;

  string report_id = "";

  //  Group: Functions
  function void build_phase(uvm_phase phase);
    string report = $sformatf("%s.build_phase", report_id);
    super.build_phase(phase);
    `uvm_info(report, $sformatf("Starting build_phase for %s", get_full_name()), UVM_NONE)

    if (!uvm_config_db#(vif_t)::get(this, "", "vif", vif))
      `uvm_fatal(report, $sformatf("Error to get vif for %s", get_full_name()))

    if (!uvm_config_db#(axis_config)::get(this, "", "m_cfg", m_cfg))
      `uvm_fatal(report, $sformatf("Error to get axis_config for %s", get_full_name()))

    transfer_ap = new("transfer_ap", this);

    `uvm_info(report, $sformatf("Finishing build_phase for %s", get_full_name()), UVM_NONE)
  endfunction : build_phase


  task run_phase(uvm_phase phase);
    string report = $sformatf("%s.run_phase", report_id);
    axis_transfer item = axis_transfer::type_id::create("item");


    super.run_phase(phase);
    `uvm_info(report, $sformatf("run_phase for %s", get_full_name()), UVM_NONE);

    forever begin
      // wait for valid data
      // if (!(vif.TVALID == 1)) @(posedge vif.TVALID);
      // if (!(vif.TREADY == 1)) @(posedge vif.TREADY);
      //do @(posedge vif.ACLK); while (!(vif.TVALID && vif.TREADY));
      wait (vif.TVALID && vif.TREADY);

      @(negedge vif.ACLK);
      if (m_cfg.TDATA_ENABLE) item.tdata <= vif.TDATA;
      if (m_cfg.TKEEP_ENABLE) item.tkeep <= vif.TKEEP;
      if (m_cfg.TLAST_ENABLE) item.tlast <= vif.TLAST;
      if (m_cfg.TSTRB_ENABLE) item.tstrb <= vif.TSTRB;
      `uvm_info(report, $sformatf("MON_%s: ITEM\n%s", m_cfg.device_type.name, item.sprint()),
                UVM_FULL)

      @(posedge vif.ACLK);
      item.timestamp = $time;
      transfer_ap.write(item);
    end

    `uvm_info(report, $sformatf("run_phase for %s", get_full_name()), UVM_NONE)
  endtask : run_phase


  function new(string name = "axis_monitor", uvm_component parent);
    super.new(name, parent);
    this.report_id = name;
  endfunction : new

endclass : axis_monitor

`endif
